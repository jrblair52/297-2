module ahb_top () (

  ahb_master master_1 (
    .host_read_1	(host_read),
    .host_write_1	(host_write),
    .host_cont_1	(host_cont),
    .host_size_1	(host_size),
    .host_addr_1	(host_addr),
    .host_wdata_1	(host_wdata),
    .bus_rdata_1	(bus_rdata),
    .bus_rdone_1	(bus_rdone),
    .bus_wready_1	(bus_wready),
    .hreset_1		(hreset),
    .hclk_1			(hclk),
    .hreset_1		(hreset),
    .hresp_1		(hresp),
    .hgrant_1		(hgrant),
    .hrdata_1		(hrdata),
    .haddr_1		(haddr),
    .hwrite_1		(hwrite),
    .hsize_1		(hsize),
    .hburst_1		(hburst),
    .hprot_1		(hprot),
    .htrans_1		(htrans),
    .hmastlock_1	(hmastlock),
    .hbusreq_1		(hbusreq),
    .hlock_1		(hlock),
    .hwdata_1		(hwdata)
  );
  
  address_decoder decoder (
    .hclk		(hclk),
    .hreset		(hreset),
    .haddr		(haddr),
    .hsel_1		(hsel_1),
    .hsel_2		(hsel_2),
    .hsel_3		(hsel_3),
    .hsel_4		(hsel_4),
    .hsel_5		(hsel_5),
    .hsel_6		(hsel_6),
    .hsel_7		(hsel_7),
    .hsel_8		(hsel_8),
    .hsel_9		(hsel_9),
    .hsel_10		(hsel_10)
    .hsel_11		(hsel_11),
    .hsel_12		(hsel_12),
    .hsel_13		(hsel_13),
    .hsel_14		(hsel_14),
    .hsel_15		(hsel_15),
    .hsel_16		(hsel_16)
  );
    
  multiplexer multiplexer (
    .haddr		(haddr),
    .hrdata_1		(hrdata_1),
    .hrdata_2		(hrdata_2),
    .hrdata_3		(hrdata_3),
    .hrdata_4		(hrdata_4),
    .hrdata_5		(hrdata_5),
    .hrdata_6		(hrdata_6),
    .hrdata_7		(hrdata_7),
    .hrdata_8		(hrdata_8),
    .hrdata_9		(hrdata_9),
    .hrdata_10		(hrdata_10),
    .hrdata_11		(hrdata_11),
    .hrdata_12		(hrdata_12),
    .hrdata_13		(hrdata_13),
    .hrdata_14		(hrdata_14),
    .hrdata_15		(hrdata_15),
    .hrdata_16		(hrdata_16),
    .hreadyout_1	(hreadyout_1),
    .hreadyout_2	(hreadyout_2),
    .hreadyout_3	(hreadyout_3),
    .hreadyout_4	(hreadyout_4),
    .hreadyout_5	(hreadyout_5),
    .hreadyout_6	(hreadyout_6),
    .hreadyout_7	(hreadyout_7),
    .hreadyout_8	(hreadyout_8),
    .hreadyout_9	(hreadyout_9),
    .hreadyout_10	(hreadyout_10),
    .hreadyout_11	(hreadyout_11),
    .hreadyout_12	(hreadyout_12),
    .hreadyout_13	(hreadyout_13),
    .hreadyout_14	(hreadyout_14),
    .hreadyout_15	(hreadyout_15),
    .hreadyout_16	(hreadyout_16),
    .hresp_1		(hresp_1),
    .hresp_2		(hresp_2),
    .hresp_3		(hresp_3),
    .hresp_4		(hresp_4),
    .hresp_5		(hresp_5),
    .hresp_6		(hresp_6),
    .hresp_7		(hresp_7),
    .hresp_8		(hresp_8),
    .hresp_9		(hresp_9),
    .hresp_10		(hresp_10),
    .hresp_11		(hresp_11),
    .hresp_12		(hresp_12),
    .hresp_13		(hresp_13),
    .hresp_14		(hresp_14),
    .hresp_15		(hresp_15),
    .hresp_16		(hresp_16),
    .hrdata		(hrdata),
    .hready		(hready),
    .hresp		(hresp)
  );
  
  ahb_arbiter arbiter (
    .hreset_n		(hreset_n),
    .hclk		(hclk),
    .hlock_0		(hlock_0),
    .hlock_1		(hlock_1),
    .hlock_2		(hlock_2),
    .hlock_3		(hlock_3),
    .hbusreq_0		(hbusreq_0),
    .hbusreq_1		(hbusreq_1),
    .hbusreq_2		(hbusreq_2),
    .hbusreq_3		(hbusreq_3),
    .addr		(haddr),
    .hsplit_0		(hsplit_0),
    .hsplit_1		(hsplit_1),
    .hsplit_2		(hsplit_2),
    .hsplit_3		(hsplit_3),
    .hburst_0		(hburst_0),
    .hresp_0		(hresp_0),
    .htrans_0		(htrans_0),
    .hready_0		(hready_0),
    .hburst_1		(hburst_1),
    .hresp_1		(hresp_1),
    .htrans_1		(htrans_1),
    .hready_1		(hready_1),
    .hburst_2		(hburst_2),
    .hresp_2		(hresp_2),
    .htrans_2		(htrans_2),
    .hready_2		(hready_2),
    .hburst_3		(hburst_3),
    .hresp_3		(hresp_3),
    .htrans_3		(htrans_3),
    .hready_3		(hready_3),
    .hgrant_1		(hgrant_1),
    .hgrant_2		(hgrant_2),
    .hgrant_3		(hgrant_3),
    .hmaster		(hmaster),
    .hmastlock		(hmastlock)
  );
  
  ahb_slave slave_1 (
    .hsel_1		(hsel),
    .hrdata_1		(hrdata)
  );
    
endmodule
